`ifndef _CONSTANT_DEFS
`define _CONSTANT_DEFS

// data bus width
`define W_DATA 32
// instruction size
`define W_INST 32
// memory address width (same for data/inst)
`define W_ADDR 32
// register file size, including 0 register
`define RF_SIZE 32
// register file address width
`define W_RFADDR 5
`define W_JADDR 26


`endif